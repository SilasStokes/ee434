* SPICE NETLIST
***************************************

.SUBCKT MUX2_X1 S A B VDD VSS Y
** N=11 EP=6 IP=0 FDC=12
M0 VSS S 1 VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=7.13e-14 AS=5.52e-14 PD=1.08e-06 PS=9.4e-07 $X=-2055 $Y=-2040 $D=1
M1 10 1 VSS VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=3.335e-14 AS=7.13e-14 PD=7.5e-07 PS=1.08e-06 $X=-1605 $Y=-2040 $D=1
M2 4 A 10 VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=7.475e-14 AS=3.335e-14 PD=1.11e-06 PS=7.5e-07 $X=-1320 $Y=-2040 $D=1
M3 11 S 4 VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=3.45e-14 AS=7.475e-14 PD=7.6e-07 PS=1.11e-06 $X=-855 $Y=-2040 $D=1
M4 VSS B 11 VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=4.715e-14 AS=3.45e-14 PD=8.7e-07 PS=7.6e-07 $X=-565 $Y=-2040 $D=1
M5 Y 4 VSS VSS NMOS_HP L=1.4e-07 W=2.3e-07 AD=4.83e-14 AS=5.75e-14 PD=8.8e-07 PS=9.6e-07 $X=210 $Y=-2030 $D=1
M6 VDD S 1 VDD PMOS_HP L=1.4e-07 W=4.05e-07 AD=1.2555e-13 AS=9.72e-14 PD=1.43e-06 PS=1.29e-06 $X=-2055 $Y=1340 $D=0
M7 6 1 VDD VDD PMOS_HP L=1.4e-07 W=4.05e-07 AD=1.39725e-13 AS=1.2555e-13 PD=1.5e-06 PS=1.43e-06 $X=-1605 $Y=1340 $D=0
M8 4 S 6 VDD PMOS_HP L=1.4e-07 W=4.05e-07 AD=9.5175e-14 AS=1.39725e-13 PD=1.28e-06 PS=1.5e-06 $X=-1120 $Y=1340 $D=0
M9 6 B 4 VDD PMOS_HP L=1.4e-07 W=4.05e-07 AD=1.3365e-13 AS=9.5175e-14 PD=1.47e-06 PS=1.28e-06 $X=-745 $Y=1340 $D=0
M10 VDD A 6 VDD PMOS_HP L=1.4e-07 W=4.05e-07 AD=1.08725e-13 AS=1.3365e-13 PD=1.5e-06 PS=1.47e-06 $X=-275 $Y=1340 $D=0
M11 Y 4 VDD VDD PMOS_HP L=1.4e-07 W=2.5e-07 AD=6.625e-14 AS=1.08725e-13 PD=1.03e-06 PS=1.5e-06 $X=210 $Y=1495 $D=0
.ENDS
***************************************
